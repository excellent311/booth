library verilog;
use verilog.vl_types.all;
entity test_mult is
end test_mult;
