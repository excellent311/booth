library verilog;
use verilog.vl_types.all;
entity bit16_cla is
    port(
        ain             : in     vl_logic_vector(15 downto 0);
        bin             : in     vl_logic_vector(15 downto 0);
        cin             : in     vl_logic;
        sum             : out    vl_logic_vector(15 downto 0);
        cout            : out    vl_logic
    );
end bit16_cla;
