library verilog;
use verilog.vl_types.all;
entity bit4_cla is
    port(
        ain             : in     vl_logic_vector(3 downto 0);
        bin             : in     vl_logic_vector(3 downto 0);
        cin             : in     vl_logic;
        sum             : out    vl_logic_vector(3 downto 0);
        cout            : out    vl_logic;
        cas_p           : out    vl_logic;
        cas_g           : out    vl_logic
    );
end bit4_cla;
