library verilog;
use verilog.vl_types.all;
entity bit4cla_logic is
    port(
        cin             : in     vl_logic;
        p3              : in     vl_logic;
        g3              : in     vl_logic;
        p2              : in     vl_logic;
        g2              : in     vl_logic;
        p1              : in     vl_logic;
        g1              : in     vl_logic;
        p0              : in     vl_logic;
        g0              : in     vl_logic;
        c3              : out    vl_logic;
        c2              : out    vl_logic;
        c1              : out    vl_logic;
        c0              : out    vl_logic
    );
end bit4cla_logic;
